module CLB (
    clk,
    A,
    B,
    C,
    D
);
  input logic clk;
  input logic A;
  input logic B;
  input logic C;
  input logic D;


endmodule
